`define ADDR_WIDTH 32
`define SIZE 2
`define BURST_SIZE 2
`define WDATA_WIDTH 32
`define RESPONSE_WIDTH 2