`define ADDR_WIDTH 32
`define DATA_WIDTH 32
`define RESPONSE_WIDTH 2
`define OUTPUT_ADDR_WIDTH 24
`define RDATA_WIDTH 32
